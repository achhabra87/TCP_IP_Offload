library verilog;
use verilog.vl_types.all;
entity pcapparser_10gbmac_test is
end pcapparser_10gbmac_test;
